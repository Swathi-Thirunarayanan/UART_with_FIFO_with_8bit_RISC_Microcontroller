----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/23/2018 02:53:40 AM
-- Design Name: 
-- Module Name: IR - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity IR is
--  Port ( );
port(
     Irin: in std_logic_vector(7 downto 0);
     clk : in std_logic;
     irload: in std_logic;
     Irout: out std_logic_vector(7 downto 0));
end IR;

architecture Behavioral of IR is

begin
process(clk,irload)
begin
if (rising_edge(clk) and (irload = '1')) then
irout <= irin;
end if;
end process;
end Behavioral;
