----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 03/23/2018 03:07:42 AM
-- Design Name: 
-- Module Name: PC - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity PC is
--  Port ( );
port(
     pcin: in std_logic_vector(7 downto 0);
     clk : in std_logic;
     rst : in std_logic;
     pcload: in std_logic;
     pcout: out std_logic_vector(7 downto 0));
end PC;

architecture Behavioral of PC is

begin

process(clk,rst,pcload)
begin
if(rst = '1') then
pcout <= x"00";
elsif (rising_edge(clk) and pcload = '1') then
pcout <= pcin;
end if;
end process;
end Behavioral;
